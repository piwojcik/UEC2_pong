/**
 * Copyright (C) 2023  AGH University of Science and Technology
 * MTM UEC2
 * Author: Piotr Kaczmarczyk
 *
 * Description:
 * Draw background.
 */


`timescale 1 ns / 1 ps

module draw_bg (
    input  logic clk,
    input  logic rst,

     vga_intf.in bg_in,
     vga_intf.out bg_out
     
);

import vga_pkg::*;


/**
 * Local variables and signals
 */

logic [11:0] rgb_nxt;


/**
 * Internal logic
 */

always_ff @(posedge clk) begin : bg_ff_blk
    if (rst) begin
        bg_out.vcount <= '0;
        bg_out.vsync  <= '0;
        bg_out.vblnk  <= '0;
        bg_out.hcount <= '0;
        bg_out.hsync  <= '0;
        bg_out.hblnk  <= '0;
        bg_out.rgb    <= '0;
    end else begin
        bg_out.vcount <= bg_in.vcount;
        bg_out.vsync  <= bg_in.vsync;
        bg_out.vblnk  <= bg_in.vblnk;
        bg_out.hcount <= bg_in.hcount;
        bg_out.hsync  <= bg_in.hsync;
        bg_out.hblnk  <= bg_in.hblnk;
        bg_out.rgb   <= rgb_nxt;
    end
end

always_comb begin : bg_comb_blk
    if (bg_in.vblnk || bg_in.hblnk) begin             // Blanking region:
        rgb_nxt = 12'h0_0_0;                   // - make it it black.
    end else begin                              // Active region:
        if (bg_in.vcount == 0)                     // - top edge:
            rgb_nxt = 12'hf_f_0;                // - - make a yellow line.
        else if (bg_in.vcount == VER_PIXELS - 1)   // - bottom edge:
            rgb_nxt = 12'hf_0_0;                // - - make a red line.
        else if (bg_in.hcount == 0)                // - left edge:
            rgb_nxt = 12'h0_f_0;                // - - make a green line.
        else if (bg_in.hcount == HOR_PIXELS - 1)   // - right edge:
            rgb_nxt = 12'h0_0_f;                // - - make a blue line.
            
        else if ((bg_in.vcount >= 25 & bg_in.vcount <= 30 & bg_in.hcount >= 100 & bg_in.hcount <= 120) |
                (bg_in.vcount >= 30 & bg_in.vcount <= 60 & bg_in.hcount >= 108 & bg_in.hcount <= 112) | 
                (bg_in.vcount >=61 & bg_in.vcount <= 65 & bg_in.hcount >= 94 & bg_in.hcount <= 108) |
                (bg_in.vcount >= 56 & bg_in.vcount <= 60 & bg_in.hcount >= 87 & bg_in.hcount <= 93))  
            rgb_nxt = 12'h1_4_f; 
        else if ((bg_in.vcount >= 25 & bg_in.vcount <= 30 & bg_in.hcount >= 145 & bg_in.hcount <= 165) |
                (bg_in.vcount >= 30 & bg_in.vcount <= 60 & bg_in.hcount >= 153 & bg_in.hcount <= 157) | 
                (bg_in.vcount >=61 & bg_in.vcount <= 65 & bg_in.hcount >= 137 & bg_in.hcount <= 153) |
                (bg_in.vcount >= 56 & bg_in.vcount <= 60 & bg_in.hcount >= 130 & bg_in.hcount <= 136))  
            rgb_nxt = 12'h1_4_f; 

        else                                    // The rest of active display pixels:
            rgb_nxt = 12'h8_8_8;                // - fill with gray.
    end
end

endmodule
